library verilog;
use verilog.vl_types.all;
entity Q6_vlg_vec_tst is
end Q6_vlg_vec_tst;
