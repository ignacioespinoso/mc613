library verilog;
use verilog.vl_types.all;
entity Q5_vlg_check_tst is
    port(
        Q5              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Q5_vlg_check_tst;
