library verilog;
use verilog.vl_types.all;
entity Q6 is
    port(
        B               : in     vl_logic;
        clk             : in     vl_logic;
        Q6              : out    vl_logic
    );
end Q6;
