library verilog;
use verilog.vl_types.all;
entity Q1_vlg_check_tst is
    port(
        Q1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Q1_vlg_check_tst;
