library verilog;
use verilog.vl_types.all;
entity Q6_vlg_check_tst is
    port(
        Q6              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Q6_vlg_check_tst;
