library verilog;
use verilog.vl_types.all;
entity Q2_vlg_check_tst is
    port(
        Q2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Q2_vlg_check_tst;
