library verilog;
use verilog.vl_types.all;
entity Maquina1_vlg_check_tst is
    port(
        z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Maquina1_vlg_check_tst;
