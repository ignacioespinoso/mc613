library verilog;
use verilog.vl_types.all;
entity Q1 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        Q1              : out    vl_logic
    );
end Q1;
