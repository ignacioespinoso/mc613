library verilog;
use verilog.vl_types.all;
entity Q3 is
    port(
        A               : in     vl_logic;
        clk             : in     vl_logic;
        Q3              : out    vl_logic
    );
end Q3;
