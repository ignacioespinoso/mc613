library verilog;
use verilog.vl_types.all;
entity Q3_vlg_vec_tst is
end Q3_vlg_vec_tst;
