library verilog;
use verilog.vl_types.all;
entity Q1_vlg_vec_tst is
end Q1_vlg_vec_tst;
