library verilog;
use verilog.vl_types.all;
entity Q5_vlg_vec_tst is
end Q5_vlg_vec_tst;
