library verilog;
use verilog.vl_types.all;
entity Q5 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        clk             : in     vl_logic;
        m               : in     vl_logic;
        n               : in     vl_logic;
        Q5              : out    vl_logic
    );
end Q5;
