library verilog;
use verilog.vl_types.all;
entity Q3_vlg_check_tst is
    port(
        Q3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Q3_vlg_check_tst;
