library verilog;
use verilog.vl_types.all;
entity Q4_vlg_check_tst is
    port(
        Q4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Q4_vlg_check_tst;
