library verilog;
use verilog.vl_types.all;
entity Q2 is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        clk             : in     vl_logic;
        Q2              : out    vl_logic
    );
end Q2;
