library verilog;
use verilog.vl_types.all;
entity Q4_vlg_vec_tst is
end Q4_vlg_vec_tst;
