library verilog;
use verilog.vl_types.all;
entity Maquina1_vlg_vec_tst is
end Maquina1_vlg_vec_tst;
