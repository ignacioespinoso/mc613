library verilog;
use verilog.vl_types.all;
entity Q2_vlg_vec_tst is
end Q2_vlg_vec_tst;
